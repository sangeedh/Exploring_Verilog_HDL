module StructuralModeling(input a, b, output c);
  and gate1(c, a, b);
endmodule
//This Verilog code demonstrates structural modeling using gate-level primitives. 
//It describes a 2-input AND gate (gate1) that connects inputs a and b to output c.
