module HelloWorld;
  initial begin
    $display("Hello, World!");
    $finish;
  end
endmodule
//This simple Verilog code prints "Hello, World!" to the console using the $display system function.
